* CMOS inverter transient test (self-contained)

.param VDD=1.8

VDD vdd 0 {VDD}
VIN in  0 PULSE(0 {VDD} 0 20p 20p 5n 10n)

MP out in vdd vdd PMOS L=180n W=1u
MN out in 0   0   NMOS L=180n W=500n

CLOAD out 0 5f

.model NMOS NMOS LEVEL=1 VTO=0.45 KP=200u LAMBDA=0.05
.model PMOS PMOS LEVEL=1 VTO=-0.45 KP=80u  LAMBDA=0.05

.tran 50p 50n

.control
  wrdata inv.csv time v(in) v(out)
.endc

.end
