* Simple CMOS Inverter
* For testing Circuit Visualization

* Power supply
VDD vdd gnd DC 1.8

* Input voltage source (can be controlled interactively)
VIN in gnd DC 0

* PMOS transistor (pulls output high when input is low)
* Format: Mdrain gate source body model W=width L=length
MP1 out in vdd vdd PMOS W=2u L=0.18u

* NMOS transistor (pulls output low when input is high)
MN1 out in gnd gnd NMOS W=1u L=0.18u

* Simple transistor models
.model NMOS NMOS (VTO=0.4 KP=200u)
.model PMOS PMOS (VTO=-0.4 KP=100u)

* DC sweep: vary input from 0 to 1.8V
.dc VIN 0 1.8 0.01

.end
