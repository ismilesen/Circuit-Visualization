* 3-stage ring oscillator using idealized behavioral inverters

.param VDD=1.8
.param VMID=0.9
.param GAIN=40

.subckt INV in out
Bdrv ndrv 0 v = { VDD * (0.5 - 0.5*tanh(GAIN*(v(in)-VMID))) }
Rout ndrv out 1k
Cout out 0 20f
.ends INV

X1 n3 n1 INV
X2 n1 n2 INV
X3 n2 n3 INV

* Break symmetry to ensure startup
.ic v(n1)=0 v(n2)=1.8 v(n3)=0

.tran 2p 20n

.control
  wrdata ring_osc_3stage.csv time v(n1) v(n2) v(n3)
.endc

.end
